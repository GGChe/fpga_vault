// Module for Hello World

module hello_word;
initial begin
    $display ("Hello World!");
    $finish;
end

endmodule //hello_word

